library work;
use work.my_package.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

entity tb is
    port (
        clk : in std_logic;
        --wink : out std_logic;
		sw_call : out std_logic;
		EEM_columns : out integer range 0 to 21 := 0;
		EEM_rows : out integer range 0 to 20 := 0;
		EEM_data: out std_logic_vector(1 to 420) := (others => '0')
    );
end entity;

architecture arch_t of tb is
	component main is
		generic(m : in integer range 0 to 6 := 6;					--metabolites
	        q : in integer range 0 to 15 := 15;					--reactions not splitted
	        qsplit : in integer range 0 to 20 := 20 ;			--reactions splitted = q + revs
	        R_rows : in integer range 0 to 20 := 20;			--qsplit
	        R_columns : in integer range 0 to 14 := 14;			--qsplit-m
	        R1_rows : in integer range 0 to 14 := 14;			--qsplit-m
			R2_rows : in integer range 0 to 6 := 6;			--m
			max_column : in integer range 0 to 100 := 100);	--max of columns in R after adding combination
	port(clock, reset : in std_logic;
	    R1_data : in std_logic_vector(1 to 196);
	    R2_data_postfix : in std_vec_array(1 to 84);
	    SW_call : out std_logic := '0';
	    EM_columns : out integer range 0 to 21 := 0;
	    EM_rows : out integer range 0 to R_rows := 0;
	    EM_data: out std_logic_vector(1 to 420) := (others => '0')
    );
	end component main;

    signal rst : std_logic := '0';
	signal RR1_data : std_logic_vector(1 to 196);
	signal RR2_data : std_vec_array(1 to 84); 
	
begin 
	
	rst <= '0';
	RR1_data <=(
		'1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0',  
		'0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
		'0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0',
		'0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1'
	);
	RR2_data <= (
		"00010000",
"00010000",
"00010000",
"00010000",
"00010000",
"11110000",
"00000000",
"00010000",
"00000000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"11110000",
"00010000",
"00000000",
"00010000",
"11110000",
"00000000",
"00010000",
"00000000",
"00000000",
"00000000",
"00010000",
"00000000",
"00000000",
"00000000",
"00010000",
"11110000",
"00000000",
"11110000",
"00010000",
"00000000",
"11110000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000",
"00100000",
"00000000",
"00000000",
"11110000",
"00010000",
"00000000",
"00010000",
"00010000",
"00000000",
"00000000",
"00000000",
"00010000",
"00000000",
"00010000",
"00000000",
"00010000",
"00010000",
"00010000",
"11110000",
"00000000",
"00010000",
"00000000",
"00000000",
"00010000",
"00000000",
"00000000",
"00000000",
"00010000",
"00000000",
"00010000",
"00000000",
"00010000",
"11110000",
"00000000",
"00010000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00010000"

	);
    --RR2_data <= ("00000000000100000000000000", "11111111111100000000000000", "11111111111100000000000000", "00000000001000000000000000", "00000000000100000000000000", "00000000000100000000000000", "11111111111100000000000000", "00000000000000000000000000");
	      
	--wink <= '1';
	
	main_comp : main generic map (6, 15, 20, 20, 14, 14, 6, 100)
					 port map (clk, rst, RR1_data, RR2_data, sw_call, EEM_columns, EEM_rows, EEM_data);
end architecture arch_t;
